../test1/dut.sv