../test1/tb_vif.sv