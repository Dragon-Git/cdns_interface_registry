../test1/testbench_pkg.sv